`define IDLE                  4'b0000
`define CHECK_TAG             4'b0001
`define WAIT_DRAM_READY       4'b0010
`define DRAM_READ             4'b0011
`define SETTLE                4'b0100
`define GIVE_TO_CPU           4'b0101
`define WAIT_DRAM_FLUSH_BLOCK 4'b0110
`define DRAM_WRITE            4'b0111
