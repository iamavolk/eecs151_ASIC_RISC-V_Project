/scratch/cs199-aly/eecs151_ASIC_RISC-V_Project/skel/build/tech-sky130-cache/sky130_ef_io.lef